�4<m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	 	 	 	 	 	 	 	 	 	 	 	                              	 	  	 	 	  	   	 	           
                   	 	   	   	  	 	 	              
               	 	  	  	  	 	  	 	                              	 	  	 	 	  	   	 	                             	 	 	 	 	 	 	 	 	 	 	 	                             	   	 	    	   	                             	  	  	  	  	  	 	                             	  	  	  	  	 	  	                           	   	 	    	   	                            	 	 	 	 	 	 	 	 	 	 	 	                                                                                                           