�4<m 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	         	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	         	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	   	 	 	 	 	 	   	      	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	           	 	      	 	 	 	 	 	 	 	 	 	 	 	 	 	 	    	 	  	 	   	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	 	 	         	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	 	 	         	 	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	 	 	       	 	 	 	 	 	      	 	 	 	 	 	 	 	 	 	                 	      	 	 	 	 	 	 	                         	 	 	 	 	 	 	             	             	 	 	 	 	 	              	            	 	 	 	 	 	 	             	  	          	 	 	 	 	 	 	      	       	    	      	 	 	 	 	 	 	 	 	 	      	    	 	 	      	 	 	   	 	 	 	 	 	 	 	 	 	      	 	 	             	 	 	 	 	 	 	 	 	 	 	 	 	      	 	             	 	 	 	 	 	 	 	 	 	 	 	 	      	 	             	 	 	 	 	 	 	 	 	 	 	 	 	 	      	             	 	 	 	 	 	 	 	 	 	 	 	 	 	 	                  	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	              	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	       	 	 	 	 	       	 	 	 	 	 	 	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	 	      	 	 	 	 	 	 	      	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 