���                                                                                                     	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	   	 	       	 	 	 	 	 	 	 	 	 	 	 	     	   	 	     	       	    	    	 	 	          	     	        
    
    	 	           	   	 	           
     	 	           	 	 	 	 	           
     	 	 	         	 	 	 	 	 	        
 
  
    
  	 	  	 	    	 	 	 	 	 	 	 	       
     
 
 
   	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	            
     	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	                 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	                	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	               	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	       	 	 	   	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	       	 	 	   	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	       	 	 	   	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	       	 	 	   	 	 	 	 	 	 	 	 	 	 	 	 
 	 	 
 	 	 
 	 	            	 	 	 	 	 	 	 	 	 	 	 
 	 	 	 
 	 	 
 	 	              	 	 	 	 	 	 	 	 	 
 	 	 
 	 	 
 	 	 
                  	 	 	 	 
 	 	 
 
   
   
                      
 	 
  
  
 
  
                       
  
  
 
  
  
                       
  
   
    
                         
   
   
                                                                                                                                                                                                      