���  	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	                                       	 	 	 	 	 	 	 	 	 	 	 	 	                                  	 	 	 	 	 	 	 	 	 	 	 	 	                                       	 	 	 	 	 	 	 	 	 	 	 	 	                                   	 	 	 	 	 	 	 	 	 	 	 	 	                                       	 	 	 	 	 	 	 	 	 	 	 	 	                               	 	 	 	 	 	 	 	 	 	 	 	 	                                       	 	 	 	 	 	 	 	 	 	 	 	 	                                  	 	 	 	 	 	 	 	 	 	 	 	 	                                       	 	 	 	 	 	 	 	 	 	 	 	 	                               	 	 	 	 	 	 	 	 	 	 	 	 	                                       	 	 	 	 	 	 	 	 	 	 	 	 	                             	 	 	 	 	 	 	 	 	 	 	 	 	                                                             	 	                                                 	 	                                                             	 	                                      	 	                                                 	 	                       	                	 	                              	                    	 	 	 	 	 	 	 	 	 	 	 	 	 	                     	 	 	 	 	 	 	 	 	 	 	 	 	 	                           	 	 	 	 	 	 	 	 	 	 	 	 	 	                     	 	 	 	 	 	 	 	 	 	 	 	 	 	                            	 	 	 	 	 	 	 	 	 	 	 	 	 	                     	 	 	 	 	 	 	 	 	 	 	 	 	 	                           	 	 	 	 	 	 	 	 	 	 	 	 	 	                     	 	 	 	 	 	 	 	 	 	 	 	 	 	                     	 	 	 	 	 	 	 	 	 	 	 	 	 	                     	 	 	 	 	 	 	 	 	 	 	 	 	 	                     	 	 	 	 	 	 	 	 	 	 	 	 	 	                                     	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	 