�4<m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 	 	 	 	 	 	 	 	 	 	 	                                	 	   	   	   	 	                         	 	      	  	 	 	                             	 	  	  	  	 	  	 	                                	 	  	 	 	  	   	 	                        	 	 	 	 	 	 	 	 	 	 	 	                                    	   	 	    	   	                        	  	  	  	  	  	 	                        	  	  	  	  	 	  	                        	   	 	    	   	                        	 	 	 	 	 	 	 	 	 	 	 	                                                                                                 