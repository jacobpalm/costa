���                                                                            
 
 
 
 
 
 
 
 
 
 
                    
 
 
 
 
 
 
   
 
 
 
 
 
                 
 
 
 
 
 
 
 
    
 
 
 
 
 
 
              
 
 
 
 
 
 
 
 
     
 
 
 
 
 
 
             
 
 
 
 
 
 
 
 
      
 
 
 
 
 
 
           
 
 
 
 
 
 
 
 
 
       
 
 
 
 
 
 
          
 
 
 
 
 
 
 
 
 
        
 
 
 
 
 
         
 
 
 
 
 
 
 
 
 
 
       
 
 
 
 
 
 
 
        
 
 
 
 
 
 
 
 
 
 
      
 
 
 
 
 
 
 
 
 
       
 
 
 
 
 
 
 
 
 
 
     
 
 
 
 
 
 
 
 
 
 
      
 
 
 
 
 
 
 
 
 
 
 
    
 
 
 
 
 
 
 
 
 
 
 
      
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
    
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
    
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
    
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
    
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
    
 
 
 
 
 
 
 
 
 
 
 
 
   
 
 
 
 
 
 
 
 
 
 
 
 
 
    
 
 
 
 
 
 
 
 
 
 
 
     
 
 
 
 
 
 
 
 
 
 
 
     
 
 
 
   
 
 
 
 
       
 
 
 
 
 
 
 
 
 
 
     
 
 
     
 
 
         
 
 
 
 
 
 
 
 
 
     
 
 
     
 
 
         
 
 
 
 
 
 
 
 
       
 
 
   
 
 
 
 
       
 
 
 
 
 
 
 
 
 
       
 
 
 
 
 
 
 
 
 
 
     
 
 
 
 
 
 
 
 
 
        
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
           
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
                   
 
 
 
 
 
 
 
 
 
 
                                            