�4<m                                                                                    	 	 	 	 	 	 	 	 	 	 	 	                       	 	   	   	   	 	                       	 	      	  	 	 	                       	 	  	  	  	 	  	 	                       	 	  	 	 	  	   	 	                         	 	 	 	 	 	 	 	 	 	 	 	                        	   	 	    	   	                        	  	  	  	  	  	 	                        	  	  	  	  	 	  	                        	   	 	    	   	                        	 	 	 	 	 	 	 	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           