�4<m         	 	 	 	 	                          	 	 	 	 	 	 	 	 	 	 	  
  
 
 
   
 
 
  
        	 	  	   	 	 	 	 	 	 	 	 
 
     
 
 
  
 
       	       	 	 	  	 	 	 	      
 
 
  
 
               	 	 	 	 	 	 	 	    
 
 
 
   
               	 	 	 	  	 	 	 	    
 
 
  
 
          	   	 	 	 	 	 	 	  	 	 	 	  
 
 
    
        	 	 	 	 	 	      	 	 	   	   
 
    
      	 	 	 	 	 	 	        	     	 
 
 
    
         	   	        	     	  
     
          	  	               	 
 
     
           	 	                 	 
 
                 	                 	 
                 	 	               	 
                  	 	              
                	 	 	                                	   	                           	 	     	 	                                   	 	                    
 
 
  
 
 
 
   	        
 
 
            
 
 
 
 
 
 
           
 
 
 
 
 
          
 
 
 
 
 
   	           
 
 
 
 
 
          
 
 
 
 
 
   	          
   
 
 
 
            
 
 
 
 
   
 	          
      
      
 
 
 
   
 
      
 	 	         
 
             
 
 
 
   
         	 	        
 
             
 
 
 
   
          	         	 	 	             
 
 
 
   
                    	 	 	            
 
 
 
   
 
 
 
 
 
                              
 
 
 
   
 
 
 
 
 
 
 
 
            
 
                
 
 
 
   
 
 
 
 
 
 
 
 
 
          
 
 
 
 
          
 
 
 
             
       
       
       
      