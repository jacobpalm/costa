�|                  ��������������   �������������y�ۜy�ۜy�ۜ��מv�lv�lv�l�ݷnonz�onz�onz��^v�onz�onz�onz��^v�v�lv�lv�l�ݷny�ۜy�ۜy�ۜ��מ�����������������������  @   @   @   �����������������y���y���y�������v��v��v���ݷ�on{�on{�on{��^w�on{�on{�on{��^w�v��v��v���ݷ�y���y���y������������������������������  @   @   @   �����������������onz�onz�onz��^v�v�lv�lv�l�ݷny�ۜy�ۜy�ۜ��מy�ۜy�ۜy�ۜ��מv�lv�lv�l�ݷnonz�onz�onz��^v��������������@   @   @   ����            �       