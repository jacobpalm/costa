���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	                                	                                	                                           
 
     
 
               
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
   
               
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
       
 
 
 
       
 
 
 
 
 
 
 
 
 
 
 
                                                                                                                                                                             