�|         0   0����000    0   0����000    ?   ?   ?����   ?   ?   ?����   0   0����    0   0����    0   0   0       0   0   0       0  ~0  ~0  ~    0  ~0  ~0  ~    ? �? �?      ? �? �?     0 �0 �0     0 �0 �0      0� ~0  ~0�     0� ~0  ~0� 
  x0�x0  0   x0�x0  0    ?��? �? `   ?��? �? ` �~0�0� 0 � �~0�0� 0 �  �0 0 �0�  �0 0 �0� ��0� `0��0 � ��0� `0��0 � ��?� ?��?  f ��?� ?��?  f ��0� `0��0 � ��0� `0��0 � ��0��0��0  ��0��0��0      