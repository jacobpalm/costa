�;y  �(br3                                                   br3                                                   brbu3urdbu3u5ld5bd6br5                                bu3u0bu2u6bd11br3                                     bu9bru2br2d2bd9br4                                    bu10ubr2dbd10br3                                      bu5bru2eu2eud2l2r6hud1gd2gd2u2l4r6br4bd7              bu7brel2r5lgeu2egr2l5regd2br4bd8br3                   bu4f2e2h4uf4uh4e2f2h2d10bd2br5                        bu4f2u10f2h2g2dfrf2d2gbd3br4                          br2bu3ueueueueul2gdglhuerbd6br4rfdglhubd5br6          bu3ue6ul5gdfreubd3frfdglhubr6bd5                      brbu3u8gdfrlgd3fr3u4rd3u3reubl2lelul3bd11br9          bu6br6g3l2hu2e4hlgdf6bd3br3                           bu10e2bd12br4                                         bu10ebd11br3                                          bu12br2g2d6fu8d8fbd2br3                               bu12br2gdgd4fdfbd2br3                                 bu2eu8fd6u6h2bd12br5                                  bu12fdfd4gdgbr5bd2                                    bu8ehfru2d4u2regfbd8br3                               bu9r2uhfregdr2l2dfhlgbd7br7                           bu7r2u2d4u2r2bd7br3                                   bu7r2u2d4u2r2bd7br2                                   bueu2ldbd3br4                                         bu1eubd3br3                                           bu7r4bd7br3                                           bu7r4bd7br3                                           bu3urdbd3br3                                          bu3 u0bd3br3                                          bu3ueueueueubd12br3                                   bu3ueueueueubd12br3                                   bu4u6ed8r3u8fd6u6hl3bd11br7                           bu5f2h2u4e2rf2d4g2lbd3br6                             bu3br2u8gerd8bd3br5                                   br3bu3u8gbd10br6                                      bu3r5l5e5ug5e5ugu2l3gbd10br8                          bu3r5l5e5u2hl2g2bd9br8                                bu4fr3u5fd3u3hl2e3lg3e3l4bd11br8                      bu4fr2e2uh2le3l5bd11br8                               br4bu3u8rd8u8lg4dr6bd6br2                             br5bu3u8g5dr6bd5br3                                   bu4fr3u5fd3u3hl4u3rd3u3r4bd11br3                      bu4fr3eu3hl4u3r5bd11br3                               bu4u5e2r2lg2d6r3u5fd3u3hl2bd8br6                      bu11br4l2g2d5fr3eu3hl3br4bd8br3                       br2bu3u3rd3u4ru4rd3u3l5br8bd11                        bu11r5dgdgdgd2br6bd3                                  bu4u2d2fr3l3u4r3l3u4gd2u2er3d8eu2bu2u2bd10br3         brbu3r3l3hu3ehuer3fdgl3r3fd3bd4br3                    bu3brr2uru7fd5u5hl3d5hu3d3fr3bd6br4                   brbu3r2e2u5hl3gd3fr4bd6br3                            bu3urdbu5uldbd8br4                                    bu3d0bu5d0bd8br3                                      bueu2ldbu5urdbd8br3                                   bueubu5d0bd8br3                                       bu7e3rg3f3lh3bd7br6                                   bu6e3g3f3bd3br3                                       bu6r5bu2l5bd8br8                                      bu4r4bu3l4br7bd7                                      bu4e3h3rf3g3bd4br5                                    bu3e3h3bd9br6                                         br2bu3urdbu3lure2ug2eu2l3gbd10br8                     br3bu3u0bu2ue3uhl3gdbd9br8                            br6bu3l4h2u3e2r4f2d2glhu2l2gdfrbd5br7                 br4bu3l2h2u3e2r3f2d2gl3huer2d3br2bd5br3               bu3u7ed8u8r3d4l3r3d4ru7bd10br3                        bu3u2r5l4u2eueudfdfd2rd2bd3br3                        bu3u8rd8r3u8l3r3d4l3r3eu2bd4d2bd4br3                  bu3u8r4fdgl3r3fd3gl3bd3br7                            bu10br5hl3d8hu6d6fr3ebd4br3                           bu10br5hl3gd6fr3ebd4br3                               bu3u8rd8r3u8fd6u6hl3br7bd11                           bu3u8r3f2d4g2l3bd3br8                                 bu3u8r4l3d4r2l2d4r3bd3br3                             bu3r4l4u4r3l3u4r4bd11br3                              bu3u8r4l3d4r2l2d4br6bd3                               bu3u4r3l3u4r4bd11br3                                  bu10br5hl3d8hu6d6fr3eu3ld3u3bd7br5                    bu7br3r2d3gl3hu6er3fbd10br3                           bu3u8rd8u4r3u4d8ru8d8bd3br3                           bu3u8d4r5u4d8bd3br3                                   bu3bru8rd8br4bd3                                      brbu3u8bd11br3                                        bu4u2rd3r3u8rd7bd4br4                                 bu5dfr3eu7bd11br3                                     bu3u8rd8u4f4rh4e4lg4bd7br8                            bu3u8d4re4g4f4bd3br3                                  bu3u8rd8r3bd3br3                                      bu3u8d8r4bd3br3                                       bu3u8f5e4ug5h4df4e5d7lu7d7bd3br4                      bu3u8f3e3d8bd3br3                                     bu3u6f6uh6uf6u6bd11br3                                bu3u8rdfdfdfdfu8bd11br3                               bu4u6ed8r3u8fd6u6hl3bd11br7                           bu4u6er3fd6gl3bd3br7                                  bu3u8rd8u4r3u4fd2u2hl3bd11br7                         bu3u8r3fd2gl3bd7br7                                   bu4u6ed8u8r3d8eu6d6gl2rfrbd2br3                       bu4u6er3fd6gl3r3hf2bd2br3                             bu3u8rd8br3u8l3r3fd2gl3r3fd3bd3br3                    bu3u8r4fd2gl4f4bd3br3                                 bu4fr2urh4uf4uh4rur2fbd10br3                          bu4fr3eu2hl3hu2er3fbd10br3                            br2bu3u8l2r5l2d8br4bd3                                bu3br3u8l3r6bd11br3                                   bu4u7rd8r3u8rd7bd4br3                                 bu11d7fr3eu7bd11br3                                   bu3u8rd8r2eu7rd6bd5br3                                bu11d2fdfdfdueueueu2bd11br3                           bu3u8rd8r3u8rd8r2eu7rd6bd5br3                         bu11d2fd2fd2u2eueudfdfd2u2eu2eu2bd11br3               bu3u3d3ru8ld3fr3u4rd3gd4ru3bd6br3                     bu3ueuehuhudfdfeueudgdgfdfdbd3br3                     bu3br2u4rd4u4l2u4ld3fr3u4rd3bd8br3                    bu11d2fdfd3u3eueu2bd11br3                             bu3r5l5u2fu2e4dg4e4u2gul4bd11br8                      bu3r4l4ueue2ueul4r4bd11br3                            bu2u10r2ld10rbd2br3                                   bu2u10rld10rbd2br3                                    bu12dfdfdfdfdbd3br3                                   bu12dfdfdfdfdbd3br3                                   bu2r2u10l2rd10bd2br4                                  bu2ru10lbd12br4                                       bu9bre2f2bd9br3                                       bu10efbd10br2                                         bu3r7bd3br2                                           bu3r7bd3br2                                           bu12f2bd10br4                                         bu11fbd10br3                                          bu8er3d6ru5d5l4u4gd2u2er4bd7br3                       bu8er2fd5l3hu2er3bd7br3                               bu3u8rd8r3u6fd4u4hl2bd9br6                            bu3u8d2r3fd4gl3bd3br4br3                              br4bu8hl2d6hu4d4fr2ebd4br3                            bu8br5hl3gd4fr3ebd4br3                                bu4u4ed6r3u8d2l2r2u2rd8bd3br3                         bu4u4er3u2d8l3r3bd3br3                                br5bu4gl3u6gd4u4er3fd2lu2d2l2bd6br6                   bu4br4gl2hu4er2fd2l3br3bd6br3                         brbu3u7gr3ld6u8r2bd11br2                              bu3bru6lr2luerbd11br3                                 bufr3u9rd8u8l4d6hu4d4fr2br5bd3                        bufr2eu8l3gd4fr3bd3br3                                bu3u8rd8u5er2d6ru5bd8br3                              bu3u8d4e2rfd5bd3br3                                   bu3u6bu2rbd2d6bd3br2                                  bu9rbu2d0bd2d6bd3br3                                  bufr2u9bu2rbd2d8bdbr3                                 brreu8lrbu2d0bd11br4                                  bu3u8rd8u2rf2rh3e3lg2bd7br6                           bu3u8d5re3g3f3bd3br3                                  bu3u8rd8bd3br3                                        bu11rd8bd3br4                                         bu3u6rd6u6r3d6ru6r3d6ru5bd8br3                        bu3u6ferfd5u4e2rfd5bd3br3                             bu3u6rd6u6r3d6ru5bd8br3                               bu3u6ferfd5bd3br3                                     bu4u4ed6r3u6l3r3fd4bd4br3                             bu4u4er2fd4gl2bd3br6                                  buu8rd8u8r3d6eu4d4gl3bd3br7                           buu8r3fd4gl3br4bd3br3                                 bu4u4ed6u6r3d6l2r2d2ru8d8bdbr3                        bu4u4er3d6l3r3d2bdbr3                                 bu3u6rd6u4e2rbd9br2                                   bu3u6fer2bd9br2                                       bu4fr2uh3uf4uh3ur2fbd8br3                             bu4fr2euhl2huer2fbd8br3                               bu4bru5lru2rd2rld6r2bd3br3                            bu11brd2lr2ld5frbd3br3                                bu4u5rd6r3u6rd6bd3br3                                 bu9d5fre2u4d6bd3br3                                   bu3u6rd6r3u6rd5bd4br3                                 bu9d2fdfdueueu2bd9br3                                 bu3u6rd6r3u6rd6r2eu5rd4bd5br3                         bu9dfdfd2u2eueudfdfd2u2eueubd9br3                     bu3u2d2ru6ld2fr3eu2ld6ru2bd5br3                       bu3ue4udg2h2udf4dbd3br3                               bufr3u3l3u6ld5fr3u6rd8bdbr3                           bufr2euhl2hu5br4d8bdbr3                               bu3r5l5e5ug5e5l5r5bd9br3                              bu9r4dg4dr4bd3br3                                     br2bu2hu3heu3ebd12br3                                 bu12br2gd3gfd3fbd2br3                                 bu2bru10bd12br4                                       bu2bru10bd12br4                                       bu2eu3ehu3hbd12br5                                    bu2eu3ehu3hbd12br5                                    bu8erfrebd9br3                                        bu10erfrebd11br3                                                                                                                                                  